library verilog;
use verilog.vl_types.all;
entity tb_filter is
end tb_filter;
