//File?tb_sram.v

`timescale 1ns/1ns

`include "sram.v"

module tb_sram();
  reg [7:0] din,addr;
  wire [7:0] dout;
  reg wr,rd,cs;
  
  sram a( dout, din, addr, wr, rd, cs );
  
  initial begin
    cs = 1'b0;
    #10 cs = 1'b1;
  end

  initial begin
    din = 8'b1010_0101;
    addr = 8'b0101_1010;
    #100 addr = 8'b1010_0101;
  end

  initial begin
    wr = 1'b0;
    rd = 1'b1;
    forever begin
        #10;
        wr = $random % 2;
        rd = $random % 2;
    end
  end

  initial begin
    $monitor("At time %4t, din=%b, addr=%b, cs=%b, wr=%b, rd=%b, dout=%b",
              $time, din, addr, cs, wr, rd, dout);
  end

endmodule
    


