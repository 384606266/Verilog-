library verilog;
use verilog.vl_types.all;
entity tb_counter8b_updown is
end tb_counter8b_updown;
