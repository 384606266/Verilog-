library verilog;
use verilog.vl_types.all;
entity tb_seq_detect is
end tb_seq_detect;
