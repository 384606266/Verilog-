library verilog;
use verilog.vl_types.all;
entity tb_shift_counter is
end tb_shift_counter;
